
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE WORK.Pack.ALL;

entity main is
	PORT (
		START : IN STD_LOGIC; -- ACTIVE HIGH
		CLK: IN STD_LOGIC;
		WRITE_BUS_DR,WRITE_BUS_AC,WRITE_BUS_IR,WRITE_BUS_MEM: inout STD_LOGIC_VECTOR(7 DOWNTO 0);
	   WRITE_BUS_AR,WRITE_BUS_PC: inout STD_LOGIC_VECTOR(7 DOWNTO 0);
		T_DEC : inout STD_LOGIC_VECTOR(2 DOWNTO 0)
		
		
		);

end main;

architecture Behavioral of main is
	-- READ_BUS : DATA FROM BUS SYSTEM TO REGISTER
	SIGNAL READ_BUS: STD_LOGIC_VECTOR(7 DOWNTO 0);
	 
	
	
	-- LOAD : TELLS REGISTER TO GET INPUT
	SIGNAL LOAD: STD_LOGIC_VECTOR(4 DOWNTO 0); --CONTROL UNIT LOAD 
	 
	-- BUS_OUT : WHEN ACTIVE, TELLS REGISTER TO OUTPUT ITS DATA
	--SIGNAL BUS_OUT: STD_LOGIC_VECTOR(7 DOWNTO 0);  --DATA FROM REGISTER TO BUS  ---------------------------------------
	
	-- _INC : CALL REGISTER INCREMENT
	SIGNAL AC_INC, PC_INC: STD_LOGIC; --CONTROL UNIT 
	
	-- CONTROL2ALU :  CONTROL UNIT OUTPUT TO  ENCODER(INPUTS) of ALU 
	SIGNAL CONTROL2ALU: STD_LOGIC_VECTOR (3 DOWNTO 0); --
	
	-- ALU_OUT
	SIGNAL ALU_OUT : STD_LOGIC_VECTOR (7 DOWNTO 0);
	
	-- COUNTER SIGNAL
	SIGNAL CLR_SQC : STD_LOGIC;
	
	-- COUNTER TO T DECODER
	--SIGNAL T_DEC : STD_LOGIC_VECTOR(2 DOWNTO 0);
	
	-- CONTROL UNIT OUTPUT HEADING TO BUS ENCODER
	SIGNAL BUS_ENC_IN : STD_LOGIC_VECTOR(7 DOWNTO 0); --INPUTS TO ENCODER OF BUS SYSTEM MUX
	
	-- BUS ENCODER OUTPUT HEADING TO COMMON BUS
	SIGNAL ENC2BUS : STD_LOGIC_VECTOR(2 DOWNTO 0); --OUTPUTS OF ENCODER OF BUS SYSTEM ( SELECT LINES OF MUX)
	
	--fixing bugs
	signal Counter_in : STD_LOGIC;
	
	-----
	--signal Data: STD_Logic_vector(7 downto 0):=(others=>'0');
	

begin
		
	-- CONNECTING REGISTERS, WIRES
	AR : REG GENERIC MAP (8) PORT MAP(READ_BUS, CLK, LOAD(0), '0', '0', '0', WRITE_BUS_AR); 
	PC : REG GENERIC MAP (8) PORT MAP(READ_BUS, CLK, LOAD(1), PC_INC, '0', START, WRITE_BUS_PC); 
	DR : REG GENERIC MAP (8) PORT MAP(READ_BUS, CLK, LOAD(2), '0', '0', '0', WRITE_BUS_DR);
	AC : REG GENERIC MAP (8) PORT MAP(ALU_OUT, CLK, LOAD(3), AC_INC, '0', '0', WRITE_BUS_AC);
	IR : REG GENERIC MAP (8) PORT MAP(READ_BUS, CLK, LOAD(4), '0', '0', '0', WRITE_BUS_IR);
	M : MEM PORT MAP(WRITE_BUS_AR(5 downto 0), WRITE_BUS_MEM, BUS_ENC_IN(6)); 

	
	 

	-- START ALU
	ALU_UNIT : ALU PORT MAP (CONTROL2ALU, WRITE_BUS_DR, WRITE_BUS_AC, ALU_OUT);
	-- END ALU 
	 
	-- COUNTERS
	Counter_in <= CLR_SQC OR START;
	T_COUNTER : COUNTER4 PORT MAP(Counter_in, CLK, '1', T_DEC);
	   
	-- CONTROL UNIT :/
	CU : CONTROL_UNIT PORT MAP (WRITE_BUS_IR(7 DOWNTO 6), T_DEC, LOAD, PC_INC, AC_INC, CLR_SQC, CONTROL2ALU, BUS_ENC_IN, WRITE_BUS_IR(1 DOWNTO 0));
  
	-- BUS ENCODER
	BUS_ENCODER : ENCODER8X3 PORT MAP (BUS_ENC_IN, ENC2BUS);
	
	-- COMMON BUS
	COMMON_BUS : COM_BUS PORT MAP (ENC2BUS, READ_BUS, WRITE_BUS_AR, WRITE_BUS_PC, WRITE_BUS_DR, WRITE_BUS_AC, WRITE_BUS_IR, WRITE_BUS_MEM);



end Behavioral; 
